library ieee;
use ieee.STD_LOGIC_1164.all;
use ieee.numeric_std.all;

entity M5_control_integral is
  port (
    clk     : in  std_logic;          -- reloj de 100 MHZ
    rst_n   : in  std_logic        -- reset del sistema (nivel bajo)
    
	-- faltan las señales por definir en el diseño de este modulo
	
	
	);  
                                                     
end entity M5_control_integral;


architecture rtl of M5_control_integral is


begin  -- architecture rtl



end architecture rtl;




